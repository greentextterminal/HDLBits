module top_module (
    output out);
    
    // creating a connection to ground
    assign out = 1'b0;
endmodule
