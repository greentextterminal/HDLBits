module top_module( 
    input a, b,
    output cout, sum 
);
    
    // Truth Table
    // a | b | s | c
    // 0 | 0 | 0 | 0
    // 0 | 1 | 1 | 0
    // 1 | 0 | 1 | 0
    // 1 | 1 | 0 | 1

    // from Truth Table the lines below can be derived
    // assign sum  = a + b;
    // assign cout = a & b;
    
    // the optimized approach is to concatenate the cout and sum and assign it with the sum of the inputs
    assign {cout, sum} = a + b;

endmodule
